module update
